-- ----------------------------------------------------------------
-- prbs.vhd
--
-- 4/8/2011 D. W. Hawkins (dwh@ovro.caltech.edu)
--
-- Pseudo-binary random sequence (PRBS) generator.
--
-- This component can be configured for a serial output or
-- parallel output. In serial output, the component is essentially
-- a linear feedback shift register (LFSR). The parallel output
-- mode can be used for transciever testing, for the generation
-- of a uniform noise source, and for the generation of Gaussian
-- noise (from the sum of uniform noise samples).
--
-- ----------------------------------------------------------------
-- Implementation description
-- --------------------------
--
-- A linear feedback shift register (LFSR) can be used to generate
-- a 1-bit PRBS. A parallel output PRBS generator generates
-- multiple PRBS bits per clock, eg. given a polynomial
-- corresponding to a PRBS7 sequence, this component can be
-- configured to generate 16-bits of the sequence every clock
-- period. The parallel output is generated by shifting the LFSR
-- state by PRBS_WIDTH effective serial clocks per clock period.
--
-- The sequence of PRBS output bits generated by an LFSR can
-- be described using a transition matrix. For example, given
-- the PRBS7 polynomial 1 + X^6 + X^7, and a Fibonacci LFSR
-- topology, the output bits can be defined in terms of the
-- transmission matrix multiplied by the 7-bit LFSR state,
-- eg., the output bit sequence for the first 20-bits of the
-- PRBS7 sequence are;
--
--      PRBS                         LFSR
--      output       0 1 2 3 4 5 6   state
--      [ p0  ] =  [ 1 0 0 0 0 0 0 ] [ s0 ]
--      [ p1  ] =  [ 0 1 0 0 0 0 0 ] [ s1 ]
--      [ p2  ] =  [ 0 0 1 0 0 0 0 ] [ s2 ]
--      [ p3  ] =  [ 0 0 0 1 0 0 0 ] [ s3 ]
--      [ p4  ] =  [ 0 0 0 0 1 0 0 ] [ s4 ]
--      [ p5  ] =  [ 0 0 0 0 0 1 0 ] [ s5 ]
--      [ p6  ] =  [ 0 0 0 0 0 0 1 ] [ s6 ]
--      [ p7  ] =  [ 1 1 0 0 0 0 0 ]
--      [ p8  ] =  [ 0 1 1 0 0 0 0 ]
--      [ p9  ] =  [ 0 0 1 1 0 0 0 ]
--      [ p10 ] =  [ 0 0 0 1 1 0 0 ]
--      [ p11 ] =  [ 0 0 0 0 1 1 0 ]
--      [ p12 ] =  [ 0 0 0 0 0 1 1 ]
--      [ p13 ] =  [ 1 1 0 0 0 0 1 ]
--      [ p14 ] =  [ 1 0 1 0 0 0 0 ]
--      [ p15 ] =  [ 0 1 0 1 0 0 0 ]
--      [ p16 ] =  [ 0 0 1 0 1 0 0 ]
--      [ p17 ] =  [ 0 0 0 1 0 1 0 ]
--      [ p18 ] =  [ 0 0 0 0 1 0 1 ]
--      [ p19 ] =  [ 1 1 0 0 0 1 0 ]
--
-- where the transition matrix consists of;
--
--  * The identity matrix in the first LFSR_WIDTH locations.
--    This is due to the fact that the first LFSR_WIDTH bits
--    in the PRBS7 sequence are the reset (or initial seed) value.
--
--  * Rows 7 and higher are constructed as the modulo-2 sum of
--    the rows 6 and 7 locations before the row, eg., the
--    row 7 value is the modulo-2 sum of row (7-6) = 1 and
--    row (7-7) = 0.
--
--    The row values can also be calculated using matrix
--    multiplies, eg. defining T as the 7x7 matrix starting
--    at p1, rows pN to pN+6 are given by T^N (matrix T
--    to the power of N). In VHDL, the calculation of row
--    sums is much simpler.
--
-- The transmission matrix determines the xor connections for
-- the output signals relative to the LFSR state, eg., the
-- value of output bit p7 is the xor of s0 and s1.
--
-- The PRBS_WIDTH generic can be 1-bit (a simple LFSR) or wider.
-- Regardless of the PRBS_WIDTH, there must be LFSR_WIDTH
-- registers to store the LFSR state. In the code below, the
-- constant DATA_WIDTH determines the internal register width
-- as the greater of LFSR_WIDTH and PRBS_WIDTH.
--
-- The parallel output PRBS is generated using using a transition
-- matrix of size 2*DATA_WIDTH x LFSR_WIDTH. The first DATA_WIDTH
-- entries are used to generate the initial 'seed' state of the
-- PRBS, while the next DATA_WIDTH entries determine the
-- 'next state' of the LFSR and PRBS outputs.
--
-- Conceptually, the LFSR_WIDTH LSBs in the 'data' register are
-- the LFSR state bits, and the remaining bits are previous
-- LFSR output (1-bit PRBS) bits stored in registers. The PRBS
-- output bits could be combinatorially generated using the
-- current LFSR state bits, but that would affect synthesis
-- timing, so registers are used (with the PRBS bits generated
-- from the previous LFSR state).
--
-- The VHDL implementation uses functions to initialize a
-- constant version of the transition matrix. The code then
-- uses the constant matrix to construct the XOR connections.
-- Since these connections are constant, this results in efficient
-- simulation and synthesis for wide PRBS output buses, eg., a
-- PRBS7 with 128-bit output generates the whole 127-bit PRBS
-- sequence plus 1-bit each clock period.
--
-- ----------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library control;
use control.utilities_pkg.all;
use control.lfsr_pkg.all;

-------------------------------------------------------------------

entity prbs is
    generic (
		-- LFSR width
        LFSR_WIDTH : integer := 7;

		-- Generator polynomial
        POLYNOMIAL : std_logic_vector := lfsr_polynomial(7);

		-- PRBS parallel output bits per clock
        PRBS_WIDTH : integer := 16
    );
    port (
        -- Clock and reset
        clk    : in  std_logic;
        rstN   : in  std_logic;

        -- Load a starting seed
        load   : in  std_logic;
        seed   : in  std_logic_vector(LFSR_WIDTH-1 downto 0);

        -- Enable control
        enable : in  std_logic;

        -- LFSR state
        lfsr_q : out std_logic_vector(LFSR_WIDTH-1 downto 0);

        -- PRBS output
        prbs_q : out std_logic_vector(PRBS_WIDTH-1 downto 0)
    );
end entity;

-------------------------------------------------------------------

architecture behave of prbs is

    -- ------------------------------------------------------------
    -- Constants
    -- ------------------------------------------------------------
    --
    -- LFSR/PRBS register width
	constant DATA_WIDTH : integer := max(LFSR_WIDTH,PRBS_WIDTH);

    -- ------------------------------------------------------------
    -- Types
    -- ------------------------------------------------------------
    --
	-- Transition matrix data type
	--
	-- * 2*DATA_WIDTH x LFSR_WIDTH
	-- * the first  DATA_WIDTH entries are used during reset
	-- * the second DATA_WIDTH entries are used to determine
	--   the next state (XOR feedback)
	--
	type prbs_matrix_t is array(0 to 2*DATA_WIDTH-1) of
		std_logic_vector(LFSR_WIDTH-1 downto 0);

    -- ------------------------------------------------------------
    -- Functions
    -- ------------------------------------------------------------
    --
	-- Transition matrix initialization
	function prbs_matrix_init return prbs_matrix_t is
		variable a : prbs_matrix_t;
	begin
		for i in 0 to 2*DATA_WIDTH-1 loop

			if (i  < LFSR_WIDTH) then

				-- Identity matrix in the first LFSR entries
				a(i)    := (others => '0');
				a(i)(i) := '1';

			else

				-- Calculate each row as the modulo-2 sum of
				-- the previous the rows with bits set in the
				-- generator polynomial, i.e., bits set in
				-- positions 1 through LFSR_WIDTH.
				--
				a(i) := (others => '0');
				for j in 1 to LFSR_WIDTH loop
					if (POLYNOMIAL(j) = '1') then
						a(i) := a(i) xor a(i-j);
					end if;
				end loop;

			end if;
		end loop;
		return a;
	end function;

	-- PRBS output bit
	--
	-- Calculate the PRBS output bit sum using the transition
	-- matrix row value (mask) and the LFSR state bits.
	--
	function prbs_sum_bit (
		mask  : std_logic_vector(LFSR_WIDTH-1 downto 0);
		state : std_logic_vector(LFSR_WIDTH-1 downto 0)) return std_logic is
		variable b : std_logic;
	begin
		-- Calculate an xor sum
		b := '0';
		for i in 0 to LFSR_WIDTH-1 loop
			if (mask(i) = '1') then
				b := b xor state(i);
			end if;
		end loop;
		return b;
	end function;

    -- ------------------------------------------------------------
    -- Signals
    -- ------------------------------------------------------------
    --
	-- PRBS/LFSR data
	signal data   : std_logic_vector(DATA_WIDTH-1 downto 0);

begin

    -- ------------------------------------------------------------
	-- PRBS/LFSR register
    -- ------------------------------------------------------------
    --
	process(clk, rstN)
		constant reset_seed :
			std_logic_vector(LFSR_WIDTH-1 downto 0) :=
				(others => '1');
		constant prbs_matrix : prbs_matrix_t := prbs_matrix_init;
	begin
		if (rstN = '0') then

			-- LFSR state bits reset to all ones
			data(LFSR_WIDTH-1 downto 0) <= reset_seed;

			-- The remaining output bits are calculated using
			-- the transition matrix (PRBS sums). The all-ones
			-- reset seed is used to determine output bits that
			-- are set or clear;
			--
			-- * output bits with an even number of xor terms
			--   get set to zero
			-- * bits with an odd number of xor terms get set
			--   to one
			--
			if (PRBS_WIDTH > LFSR_WIDTH) then
				for i in LFSR_WIDTH to PRBS_WIDTH-1 loop
					data(i)  <=
						prbs_sum_bit(prbs_matrix(i), reset_seed);
				end loop;
			end if;

		elsif rising_edge(clk) then

			if (load = '1') then
				-- LFSR state bits get loaded with seed
				data(LFSR_WIDTH-1 downto 0) <= seed;

				-- Others bits calculated based on seed
				if (PRBS_WIDTH > LFSR_WIDTH) then
					for i in LFSR_WIDTH to PRBS_WIDTH-1 loop
						data(i)  <=
							prbs_sum_bit(prbs_matrix(i), seed);
					end loop;
				end if;

			elsif (enable = '1') then

				-- PRBS parallel output update
				-- * the current LFSR state is encoded in
				--   data(LFSR_WIDTH-1 downto 0)
				-- * the next PRBS output is PRBS_WIDTH states
				--   further on from the current state.
				--
				for i in 0 to DATA_WIDTH-1 loop
					data(i)  <=
						prbs_sum_bit(prbs_matrix(i+PRBS_WIDTH),
							data(LFSR_WIDTH-1 downto 0));
				end loop;

			end if;
		end if;
	end process;

	-- LFSR state output
	lfsr_q <= data(LFSR_WIDTH-1 downto 0);

	-- PRBS parallel output
	prbs_q <= data(PRBS_WIDTH-1 downto 0);

end architecture;

